// soc_system.v

// Generated using ACDS version 21.1 842

`timescale 1 ps / 1 ps
module soc_system (
		input  wire [7:0]  apple_sprite_s1_address,                      //                  apple_sprite_s1.address
		input  wire        apple_sprite_s1_debugaccess,                  //                                 .debugaccess
		input  wire        apple_sprite_s1_clken,                        //                                 .clken
		input  wire        apple_sprite_s1_chipselect,                   //                                 .chipselect
		input  wire        apple_sprite_s1_write,                        //                                 .write
		output wire [15:0] apple_sprite_s1_readdata,                     //                                 .readdata
		input  wire [15:0] apple_sprite_s1_writedata,                    //                                 .writedata
		input  wire [1:0]  apple_sprite_s1_byteenable,                   //                                 .byteenable
		input  wire        clk_clk,                                      //                              clk.clk
		output wire        hps_hps_io_emac1_inst_TX_CLK,                 //                              hps.hps_io_emac1_inst_TX_CLK
		output wire        hps_hps_io_emac1_inst_TXD0,                   //                                 .hps_io_emac1_inst_TXD0
		output wire        hps_hps_io_emac1_inst_TXD1,                   //                                 .hps_io_emac1_inst_TXD1
		output wire        hps_hps_io_emac1_inst_TXD2,                   //                                 .hps_io_emac1_inst_TXD2
		output wire        hps_hps_io_emac1_inst_TXD3,                   //                                 .hps_io_emac1_inst_TXD3
		input  wire        hps_hps_io_emac1_inst_RXD0,                   //                                 .hps_io_emac1_inst_RXD0
		inout  wire        hps_hps_io_emac1_inst_MDIO,                   //                                 .hps_io_emac1_inst_MDIO
		output wire        hps_hps_io_emac1_inst_MDC,                    //                                 .hps_io_emac1_inst_MDC
		input  wire        hps_hps_io_emac1_inst_RX_CTL,                 //                                 .hps_io_emac1_inst_RX_CTL
		output wire        hps_hps_io_emac1_inst_TX_CTL,                 //                                 .hps_io_emac1_inst_TX_CTL
		input  wire        hps_hps_io_emac1_inst_RX_CLK,                 //                                 .hps_io_emac1_inst_RX_CLK
		input  wire        hps_hps_io_emac1_inst_RXD1,                   //                                 .hps_io_emac1_inst_RXD1
		input  wire        hps_hps_io_emac1_inst_RXD2,                   //                                 .hps_io_emac1_inst_RXD2
		input  wire        hps_hps_io_emac1_inst_RXD3,                   //                                 .hps_io_emac1_inst_RXD3
		inout  wire        hps_hps_io_sdio_inst_CMD,                     //                                 .hps_io_sdio_inst_CMD
		inout  wire        hps_hps_io_sdio_inst_D0,                      //                                 .hps_io_sdio_inst_D0
		inout  wire        hps_hps_io_sdio_inst_D1,                      //                                 .hps_io_sdio_inst_D1
		output wire        hps_hps_io_sdio_inst_CLK,                     //                                 .hps_io_sdio_inst_CLK
		inout  wire        hps_hps_io_sdio_inst_D2,                      //                                 .hps_io_sdio_inst_D2
		inout  wire        hps_hps_io_sdio_inst_D3,                      //                                 .hps_io_sdio_inst_D3
		inout  wire        hps_hps_io_usb1_inst_D0,                      //                                 .hps_io_usb1_inst_D0
		inout  wire        hps_hps_io_usb1_inst_D1,                      //                                 .hps_io_usb1_inst_D1
		inout  wire        hps_hps_io_usb1_inst_D2,                      //                                 .hps_io_usb1_inst_D2
		inout  wire        hps_hps_io_usb1_inst_D3,                      //                                 .hps_io_usb1_inst_D3
		inout  wire        hps_hps_io_usb1_inst_D4,                      //                                 .hps_io_usb1_inst_D4
		inout  wire        hps_hps_io_usb1_inst_D5,                      //                                 .hps_io_usb1_inst_D5
		inout  wire        hps_hps_io_usb1_inst_D6,                      //                                 .hps_io_usb1_inst_D6
		inout  wire        hps_hps_io_usb1_inst_D7,                      //                                 .hps_io_usb1_inst_D7
		input  wire        hps_hps_io_usb1_inst_CLK,                     //                                 .hps_io_usb1_inst_CLK
		output wire        hps_hps_io_usb1_inst_STP,                     //                                 .hps_io_usb1_inst_STP
		input  wire        hps_hps_io_usb1_inst_DIR,                     //                                 .hps_io_usb1_inst_DIR
		input  wire        hps_hps_io_usb1_inst_NXT,                     //                                 .hps_io_usb1_inst_NXT
		output wire        hps_hps_io_spim1_inst_CLK,                    //                                 .hps_io_spim1_inst_CLK
		output wire        hps_hps_io_spim1_inst_MOSI,                   //                                 .hps_io_spim1_inst_MOSI
		input  wire        hps_hps_io_spim1_inst_MISO,                   //                                 .hps_io_spim1_inst_MISO
		output wire        hps_hps_io_spim1_inst_SS0,                    //                                 .hps_io_spim1_inst_SS0
		input  wire        hps_hps_io_uart0_inst_RX,                     //                                 .hps_io_uart0_inst_RX
		output wire        hps_hps_io_uart0_inst_TX,                     //                                 .hps_io_uart0_inst_TX
		inout  wire        hps_hps_io_i2c0_inst_SDA,                     //                                 .hps_io_i2c0_inst_SDA
		inout  wire        hps_hps_io_i2c0_inst_SCL,                     //                                 .hps_io_i2c0_inst_SCL
		inout  wire        hps_hps_io_i2c1_inst_SDA,                     //                                 .hps_io_i2c1_inst_SDA
		inout  wire        hps_hps_io_i2c1_inst_SCL,                     //                                 .hps_io_i2c1_inst_SCL
		inout  wire        hps_hps_io_gpio_inst_GPIO09,                  //                                 .hps_io_gpio_inst_GPIO09
		inout  wire        hps_hps_io_gpio_inst_GPIO35,                  //                                 .hps_io_gpio_inst_GPIO35
		inout  wire        hps_hps_io_gpio_inst_GPIO40,                  //                                 .hps_io_gpio_inst_GPIO40
		inout  wire        hps_hps_io_gpio_inst_GPIO48,                  //                                 .hps_io_gpio_inst_GPIO48
		inout  wire        hps_hps_io_gpio_inst_GPIO53,                  //                                 .hps_io_gpio_inst_GPIO53
		inout  wire        hps_hps_io_gpio_inst_GPIO54,                  //                                 .hps_io_gpio_inst_GPIO54
		inout  wire        hps_hps_io_gpio_inst_GPIO61,                  //                                 .hps_io_gpio_inst_GPIO61
		output wire [14:0] hps_ddr3_mem_a,                               //                         hps_ddr3.mem_a
		output wire [2:0]  hps_ddr3_mem_ba,                              //                                 .mem_ba
		output wire        hps_ddr3_mem_ck,                              //                                 .mem_ck
		output wire        hps_ddr3_mem_ck_n,                            //                                 .mem_ck_n
		output wire        hps_ddr3_mem_cke,                             //                                 .mem_cke
		output wire        hps_ddr3_mem_cs_n,                            //                                 .mem_cs_n
		output wire        hps_ddr3_mem_ras_n,                           //                                 .mem_ras_n
		output wire        hps_ddr3_mem_cas_n,                           //                                 .mem_cas_n
		output wire        hps_ddr3_mem_we_n,                            //                                 .mem_we_n
		output wire        hps_ddr3_mem_reset_n,                         //                                 .mem_reset_n
		inout  wire [31:0] hps_ddr3_mem_dq,                              //                                 .mem_dq
		inout  wire [3:0]  hps_ddr3_mem_dqs,                             //                                 .mem_dqs
		inout  wire [3:0]  hps_ddr3_mem_dqs_n,                           //                                 .mem_dqs_n
		output wire        hps_ddr3_mem_odt,                             //                                 .mem_odt
		output wire [3:0]  hps_ddr3_mem_dm,                              //                                 .mem_dm
		input  wire        hps_ddr3_oct_rzqin,                           //                                 .oct_rzqin
		input  wire [2:0]  map1_0_avalon_slave_0_address,                //            map1_0_avalon_slave_0.address
		input  wire        map1_0_avalon_slave_0_chipselect,             //                                 .chipselect
		input  wire        map1_0_avalon_slave_0_write,                  //                                 .write
		input  wire [7:0]  map1_0_avalon_slave_0_writedata,              //                                 .writedata
		output wire [7:0]  map1_0_vga_b,                                 //                       map1_0_vga.b
		output wire        map1_0_vga_blank_n,                           //                                 .blank_n
		output wire        map1_0_vga_clk,                               //                                 .clk
		output wire [7:0]  map1_0_vga_g,                                 //                                 .g
		output wire        map1_0_vga_hs,                                //                                 .hs
		output wire [7:0]  map1_0_vga_r,                                 //                                 .r
		output wire        map1_0_vga_sync_n,                            //                                 .sync_n
		output wire        map1_0_vga_vs,                                //                                 .vs
		input  wire [2:0]  map1_1_avalon_slave_0_address,                //            map1_1_avalon_slave_0.address
		input  wire        map1_1_avalon_slave_0_chipselect,             //                                 .chipselect
		input  wire        map1_1_avalon_slave_0_write,                  //                                 .write
		input  wire [7:0]  map1_1_avalon_slave_0_writedata,              //                                 .writedata
		output wire [7:0]  map1_1_vga_b,                                 //                       map1_1_vga.b
		output wire        map1_1_vga_blank_n,                           //                                 .blank_n
		output wire        map1_1_vga_clk,                               //                                 .clk
		output wire [7:0]  map1_1_vga_g,                                 //                                 .g
		output wire        map1_1_vga_hs,                                //                                 .hs
		output wire [7:0]  map1_1_vga_r,                                 //                                 .r
		output wire        map1_1_vga_sync_n,                            //                                 .sync_n
		output wire        map1_1_vga_vs,                                //                                 .vs
		input  wire        reset_reset_n,                                //                            reset.reset_n
		input  wire [7:0]  snake_body_bottomleft_sprite_s1_address,      //  snake_body_bottomleft_sprite_s1.address
		input  wire        snake_body_bottomleft_sprite_s1_debugaccess,  //                                 .debugaccess
		input  wire        snake_body_bottomleft_sprite_s1_clken,        //                                 .clken
		input  wire        snake_body_bottomleft_sprite_s1_chipselect,   //                                 .chipselect
		input  wire        snake_body_bottomleft_sprite_s1_write,        //                                 .write
		output wire [15:0] snake_body_bottomleft_sprite_s1_readdata,     //                                 .readdata
		input  wire [15:0] snake_body_bottomleft_sprite_s1_writedata,    //                                 .writedata
		input  wire [1:0]  snake_body_bottomleft_sprite_s1_byteenable,   //                                 .byteenable
		input  wire [7:0]  snake_body_bottomright_sprite_s1_address,     // snake_body_bottomright_sprite_s1.address
		input  wire        snake_body_bottomright_sprite_s1_debugaccess, //                                 .debugaccess
		input  wire        snake_body_bottomright_sprite_s1_clken,       //                                 .clken
		input  wire        snake_body_bottomright_sprite_s1_chipselect,  //                                 .chipselect
		input  wire        snake_body_bottomright_sprite_s1_write,       //                                 .write
		output wire [15:0] snake_body_bottomright_sprite_s1_readdata,    //                                 .readdata
		input  wire [15:0] snake_body_bottomright_sprite_s1_writedata,   //                                 .writedata
		input  wire [1:0]  snake_body_bottomright_sprite_s1_byteenable,  //                                 .byteenable
		input  wire [7:0]  snake_body_horizontal_sprite_s1_address,      //  snake_body_horizontal_sprite_s1.address
		input  wire        snake_body_horizontal_sprite_s1_debugaccess,  //                                 .debugaccess
		input  wire        snake_body_horizontal_sprite_s1_clken,        //                                 .clken
		input  wire        snake_body_horizontal_sprite_s1_chipselect,   //                                 .chipselect
		input  wire        snake_body_horizontal_sprite_s1_write,        //                                 .write
		output wire [15:0] snake_body_horizontal_sprite_s1_readdata,     //                                 .readdata
		input  wire [15:0] snake_body_horizontal_sprite_s1_writedata,    //                                 .writedata
		input  wire [1:0]  snake_body_horizontal_sprite_s1_byteenable,   //                                 .byteenable
		input  wire [7:0]  snake_body_topleft_sprite_s1_address,         //     snake_body_topleft_sprite_s1.address
		input  wire        snake_body_topleft_sprite_s1_debugaccess,     //                                 .debugaccess
		input  wire        snake_body_topleft_sprite_s1_clken,           //                                 .clken
		input  wire        snake_body_topleft_sprite_s1_chipselect,      //                                 .chipselect
		input  wire        snake_body_topleft_sprite_s1_write,           //                                 .write
		output wire [15:0] snake_body_topleft_sprite_s1_readdata,        //                                 .readdata
		input  wire [15:0] snake_body_topleft_sprite_s1_writedata,       //                                 .writedata
		input  wire [1:0]  snake_body_topleft_sprite_s1_byteenable,      //                                 .byteenable
		input  wire [7:0]  snake_body_topright_sprite_s1_address,        //    snake_body_topright_sprite_s1.address
		input  wire        snake_body_topright_sprite_s1_debugaccess,    //                                 .debugaccess
		input  wire        snake_body_topright_sprite_s1_clken,          //                                 .clken
		input  wire        snake_body_topright_sprite_s1_chipselect,     //                                 .chipselect
		input  wire        snake_body_topright_sprite_s1_write,          //                                 .write
		output wire [15:0] snake_body_topright_sprite_s1_readdata,       //                                 .readdata
		input  wire [15:0] snake_body_topright_sprite_s1_writedata,      //                                 .writedata
		input  wire [1:0]  snake_body_topright_sprite_s1_byteenable,     //                                 .byteenable
		input  wire [7:0]  snake_body_vertical_sprite_s1_address,        //    snake_body_vertical_sprite_s1.address
		input  wire        snake_body_vertical_sprite_s1_debugaccess,    //                                 .debugaccess
		input  wire        snake_body_vertical_sprite_s1_clken,          //                                 .clken
		input  wire        snake_body_vertical_sprite_s1_chipselect,     //                                 .chipselect
		input  wire        snake_body_vertical_sprite_s1_write,          //                                 .write
		output wire [15:0] snake_body_vertical_sprite_s1_readdata,       //                                 .readdata
		input  wire [15:0] snake_body_vertical_sprite_s1_writedata,      //                                 .writedata
		input  wire [1:0]  snake_body_vertical_sprite_s1_byteenable,     //                                 .byteenable
		input  wire [7:0]  snake_head_down_sprite_s1_address,            //        snake_head_down_sprite_s1.address
		input  wire        snake_head_down_sprite_s1_debugaccess,        //                                 .debugaccess
		input  wire        snake_head_down_sprite_s1_clken,              //                                 .clken
		input  wire        snake_head_down_sprite_s1_chipselect,         //                                 .chipselect
		input  wire        snake_head_down_sprite_s1_write,              //                                 .write
		output wire [15:0] snake_head_down_sprite_s1_readdata,           //                                 .readdata
		input  wire [15:0] snake_head_down_sprite_s1_writedata,          //                                 .writedata
		input  wire [1:0]  snake_head_down_sprite_s1_byteenable,         //                                 .byteenable
		input  wire [7:0]  snake_head_left_sprite_s1_address,            //        snake_head_left_sprite_s1.address
		input  wire        snake_head_left_sprite_s1_debugaccess,        //                                 .debugaccess
		input  wire        snake_head_left_sprite_s1_clken,              //                                 .clken
		input  wire        snake_head_left_sprite_s1_chipselect,         //                                 .chipselect
		input  wire        snake_head_left_sprite_s1_write,              //                                 .write
		output wire [15:0] snake_head_left_sprite_s1_readdata,           //                                 .readdata
		input  wire [15:0] snake_head_left_sprite_s1_writedata,          //                                 .writedata
		input  wire [1:0]  snake_head_left_sprite_s1_byteenable,         //                                 .byteenable
		input  wire [7:0]  snake_head_right_sprite_s1_address,           //       snake_head_right_sprite_s1.address
		input  wire        snake_head_right_sprite_s1_debugaccess,       //                                 .debugaccess
		input  wire        snake_head_right_sprite_s1_clken,             //                                 .clken
		input  wire        snake_head_right_sprite_s1_chipselect,        //                                 .chipselect
		input  wire        snake_head_right_sprite_s1_write,             //                                 .write
		output wire [15:0] snake_head_right_sprite_s1_readdata,          //                                 .readdata
		input  wire [15:0] snake_head_right_sprite_s1_writedata,         //                                 .writedata
		input  wire [1:0]  snake_head_right_sprite_s1_byteenable,        //                                 .byteenable
		input  wire [7:0]  snake_head_up_sprite_s1_address,              //          snake_head_up_sprite_s1.address
		input  wire        snake_head_up_sprite_s1_debugaccess,          //                                 .debugaccess
		input  wire        snake_head_up_sprite_s1_clken,                //                                 .clken
		input  wire        snake_head_up_sprite_s1_chipselect,           //                                 .chipselect
		input  wire        snake_head_up_sprite_s1_write,                //                                 .write
		output wire [15:0] snake_head_up_sprite_s1_readdata,             //                                 .readdata
		input  wire [15:0] snake_head_up_sprite_s1_writedata,            //                                 .writedata
		input  wire [1:0]  snake_head_up_sprite_s1_byteenable,           //                                 .byteenable
		input  wire [7:0]  snake_tail_down_sprite_s1_address,            //        snake_tail_down_sprite_s1.address
		input  wire        snake_tail_down_sprite_s1_debugaccess,        //                                 .debugaccess
		input  wire        snake_tail_down_sprite_s1_clken,              //                                 .clken
		input  wire        snake_tail_down_sprite_s1_chipselect,         //                                 .chipselect
		input  wire        snake_tail_down_sprite_s1_write,              //                                 .write
		output wire [15:0] snake_tail_down_sprite_s1_readdata,           //                                 .readdata
		input  wire [15:0] snake_tail_down_sprite_s1_writedata,          //                                 .writedata
		input  wire [1:0]  snake_tail_down_sprite_s1_byteenable,         //                                 .byteenable
		input  wire [7:0]  snake_tail_left_sprite_s1_address,            //        snake_tail_left_sprite_s1.address
		input  wire        snake_tail_left_sprite_s1_debugaccess,        //                                 .debugaccess
		input  wire        snake_tail_left_sprite_s1_clken,              //                                 .clken
		input  wire        snake_tail_left_sprite_s1_chipselect,         //                                 .chipselect
		input  wire        snake_tail_left_sprite_s1_write,              //                                 .write
		output wire [15:0] snake_tail_left_sprite_s1_readdata,           //                                 .readdata
		input  wire [15:0] snake_tail_left_sprite_s1_writedata,          //                                 .writedata
		input  wire [1:0]  snake_tail_left_sprite_s1_byteenable,         //                                 .byteenable
		input  wire [7:0]  snake_tail_right_sprite_s1_address,           //       snake_tail_right_sprite_s1.address
		input  wire        snake_tail_right_sprite_s1_debugaccess,       //                                 .debugaccess
		input  wire        snake_tail_right_sprite_s1_clken,             //                                 .clken
		input  wire        snake_tail_right_sprite_s1_chipselect,        //                                 .chipselect
		input  wire        snake_tail_right_sprite_s1_write,             //                                 .write
		output wire [15:0] snake_tail_right_sprite_s1_readdata,          //                                 .readdata
		input  wire [15:0] snake_tail_right_sprite_s1_writedata,         //                                 .writedata
		input  wire [1:0]  snake_tail_right_sprite_s1_byteenable,        //                                 .byteenable
		output wire [7:0]  vga_b,                                        //                              vga.b
		output wire        vga_blank_n,                                  //                                 .blank_n
		output wire        vga_clk,                                      //                                 .clk
		output wire [7:0]  vga_g,                                        //                                 .g
		output wire        vga_hs,                                       //                                 .hs
		output wire [7:0]  vga_r,                                        //                                 .r
		output wire        vga_sync_n,                                   //                                 .sync_n
		output wire        vga_vs,                                       //                                 .vs
		input  wire [9:0]  wall_sprite_s1_address,                       //                   wall_sprite_s1.address
		input  wire        wall_sprite_s1_debugaccess,                   //                                 .debugaccess
		input  wire        wall_sprite_s1_clken,                         //                                 .clken
		input  wire        wall_sprite_s1_chipselect,                    //                                 .chipselect
		input  wire        wall_sprite_s1_write,                         //                                 .write
		output wire [15:0] wall_sprite_s1_readdata,                      //                                 .readdata
		input  wire [15:0] wall_sprite_s1_writedata,                     //                                 .writedata
		input  wire [1:0]  wall_sprite_s1_byteenable                     //                                 .byteenable
	);

	wire   [1:0] hps_0_h2f_axi_master_awburst;                           // hps_0:h2f_AWBURST -> mm_interconnect_0:hps_0_h2f_axi_master_awburst
	wire   [3:0] hps_0_h2f_axi_master_arlen;                             // hps_0:h2f_ARLEN -> mm_interconnect_0:hps_0_h2f_axi_master_arlen
	wire   [7:0] hps_0_h2f_axi_master_wstrb;                             // hps_0:h2f_WSTRB -> mm_interconnect_0:hps_0_h2f_axi_master_wstrb
	wire         hps_0_h2f_axi_master_wready;                            // mm_interconnect_0:hps_0_h2f_axi_master_wready -> hps_0:h2f_WREADY
	wire  [11:0] hps_0_h2f_axi_master_rid;                               // mm_interconnect_0:hps_0_h2f_axi_master_rid -> hps_0:h2f_RID
	wire         hps_0_h2f_axi_master_rready;                            // hps_0:h2f_RREADY -> mm_interconnect_0:hps_0_h2f_axi_master_rready
	wire   [3:0] hps_0_h2f_axi_master_awlen;                             // hps_0:h2f_AWLEN -> mm_interconnect_0:hps_0_h2f_axi_master_awlen
	wire  [11:0] hps_0_h2f_axi_master_wid;                               // hps_0:h2f_WID -> mm_interconnect_0:hps_0_h2f_axi_master_wid
	wire   [3:0] hps_0_h2f_axi_master_arcache;                           // hps_0:h2f_ARCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_arcache
	wire         hps_0_h2f_axi_master_wvalid;                            // hps_0:h2f_WVALID -> mm_interconnect_0:hps_0_h2f_axi_master_wvalid
	wire  [29:0] hps_0_h2f_axi_master_araddr;                            // hps_0:h2f_ARADDR -> mm_interconnect_0:hps_0_h2f_axi_master_araddr
	wire   [2:0] hps_0_h2f_axi_master_arprot;                            // hps_0:h2f_ARPROT -> mm_interconnect_0:hps_0_h2f_axi_master_arprot
	wire   [2:0] hps_0_h2f_axi_master_awprot;                            // hps_0:h2f_AWPROT -> mm_interconnect_0:hps_0_h2f_axi_master_awprot
	wire  [63:0] hps_0_h2f_axi_master_wdata;                             // hps_0:h2f_WDATA -> mm_interconnect_0:hps_0_h2f_axi_master_wdata
	wire         hps_0_h2f_axi_master_arvalid;                           // hps_0:h2f_ARVALID -> mm_interconnect_0:hps_0_h2f_axi_master_arvalid
	wire   [3:0] hps_0_h2f_axi_master_awcache;                           // hps_0:h2f_AWCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_awcache
	wire  [11:0] hps_0_h2f_axi_master_arid;                              // hps_0:h2f_ARID -> mm_interconnect_0:hps_0_h2f_axi_master_arid
	wire   [1:0] hps_0_h2f_axi_master_arlock;                            // hps_0:h2f_ARLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_arlock
	wire   [1:0] hps_0_h2f_axi_master_awlock;                            // hps_0:h2f_AWLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_awlock
	wire  [29:0] hps_0_h2f_axi_master_awaddr;                            // hps_0:h2f_AWADDR -> mm_interconnect_0:hps_0_h2f_axi_master_awaddr
	wire   [1:0] hps_0_h2f_axi_master_bresp;                             // mm_interconnect_0:hps_0_h2f_axi_master_bresp -> hps_0:h2f_BRESP
	wire         hps_0_h2f_axi_master_arready;                           // mm_interconnect_0:hps_0_h2f_axi_master_arready -> hps_0:h2f_ARREADY
	wire  [63:0] hps_0_h2f_axi_master_rdata;                             // mm_interconnect_0:hps_0_h2f_axi_master_rdata -> hps_0:h2f_RDATA
	wire         hps_0_h2f_axi_master_awready;                           // mm_interconnect_0:hps_0_h2f_axi_master_awready -> hps_0:h2f_AWREADY
	wire   [1:0] hps_0_h2f_axi_master_arburst;                           // hps_0:h2f_ARBURST -> mm_interconnect_0:hps_0_h2f_axi_master_arburst
	wire   [2:0] hps_0_h2f_axi_master_arsize;                            // hps_0:h2f_ARSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_arsize
	wire         hps_0_h2f_axi_master_bready;                            // hps_0:h2f_BREADY -> mm_interconnect_0:hps_0_h2f_axi_master_bready
	wire         hps_0_h2f_axi_master_rlast;                             // mm_interconnect_0:hps_0_h2f_axi_master_rlast -> hps_0:h2f_RLAST
	wire         hps_0_h2f_axi_master_wlast;                             // hps_0:h2f_WLAST -> mm_interconnect_0:hps_0_h2f_axi_master_wlast
	wire   [1:0] hps_0_h2f_axi_master_rresp;                             // mm_interconnect_0:hps_0_h2f_axi_master_rresp -> hps_0:h2f_RRESP
	wire  [11:0] hps_0_h2f_axi_master_awid;                              // hps_0:h2f_AWID -> mm_interconnect_0:hps_0_h2f_axi_master_awid
	wire  [11:0] hps_0_h2f_axi_master_bid;                               // mm_interconnect_0:hps_0_h2f_axi_master_bid -> hps_0:h2f_BID
	wire         hps_0_h2f_axi_master_bvalid;                            // mm_interconnect_0:hps_0_h2f_axi_master_bvalid -> hps_0:h2f_BVALID
	wire   [2:0] hps_0_h2f_axi_master_awsize;                            // hps_0:h2f_AWSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_awsize
	wire         hps_0_h2f_axi_master_awvalid;                           // hps_0:h2f_AWVALID -> mm_interconnect_0:hps_0_h2f_axi_master_awvalid
	wire         hps_0_h2f_axi_master_rvalid;                            // mm_interconnect_0:hps_0_h2f_axi_master_rvalid -> hps_0:h2f_RVALID
	wire         mm_interconnect_0_snake_tail_up_sprite_s1_chipselect;   // mm_interconnect_0:snake_tail_up_sprite_s1_chipselect -> snake_tail_up_sprite:chipselect
	wire  [15:0] mm_interconnect_0_snake_tail_up_sprite_s1_readdata;     // snake_tail_up_sprite:readdata -> mm_interconnect_0:snake_tail_up_sprite_s1_readdata
	wire         mm_interconnect_0_snake_tail_up_sprite_s1_debugaccess;  // mm_interconnect_0:snake_tail_up_sprite_s1_debugaccess -> snake_tail_up_sprite:debugaccess
	wire   [7:0] mm_interconnect_0_snake_tail_up_sprite_s1_address;      // mm_interconnect_0:snake_tail_up_sprite_s1_address -> snake_tail_up_sprite:address
	wire   [1:0] mm_interconnect_0_snake_tail_up_sprite_s1_byteenable;   // mm_interconnect_0:snake_tail_up_sprite_s1_byteenable -> snake_tail_up_sprite:byteenable
	wire         mm_interconnect_0_snake_tail_up_sprite_s1_write;        // mm_interconnect_0:snake_tail_up_sprite_s1_write -> snake_tail_up_sprite:write
	wire  [15:0] mm_interconnect_0_snake_tail_up_sprite_s1_writedata;    // mm_interconnect_0:snake_tail_up_sprite_s1_writedata -> snake_tail_up_sprite:writedata
	wire         mm_interconnect_0_snake_tail_up_sprite_s1_clken;        // mm_interconnect_0:snake_tail_up_sprite_s1_clken -> snake_tail_up_sprite:clken
	wire   [1:0] hps_0_h2f_lw_axi_master_awburst;                        // hps_0:h2f_lw_AWBURST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awburst
	wire   [3:0] hps_0_h2f_lw_axi_master_arlen;                          // hps_0:h2f_lw_ARLEN -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arlen
	wire   [3:0] hps_0_h2f_lw_axi_master_wstrb;                          // hps_0:h2f_lw_WSTRB -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wstrb
	wire         hps_0_h2f_lw_axi_master_wready;                         // mm_interconnect_1:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire  [11:0] hps_0_h2f_lw_axi_master_rid;                            // mm_interconnect_1:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire         hps_0_h2f_lw_axi_master_rready;                         // hps_0:h2f_lw_RREADY -> mm_interconnect_1:hps_0_h2f_lw_axi_master_rready
	wire   [3:0] hps_0_h2f_lw_axi_master_awlen;                          // hps_0:h2f_lw_AWLEN -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awlen
	wire  [11:0] hps_0_h2f_lw_axi_master_wid;                            // hps_0:h2f_lw_WID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wid
	wire   [3:0] hps_0_h2f_lw_axi_master_arcache;                        // hps_0:h2f_lw_ARCACHE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arcache
	wire         hps_0_h2f_lw_axi_master_wvalid;                         // hps_0:h2f_lw_WVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wvalid
	wire  [20:0] hps_0_h2f_lw_axi_master_araddr;                         // hps_0:h2f_lw_ARADDR -> mm_interconnect_1:hps_0_h2f_lw_axi_master_araddr
	wire   [2:0] hps_0_h2f_lw_axi_master_arprot;                         // hps_0:h2f_lw_ARPROT -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arprot
	wire   [2:0] hps_0_h2f_lw_axi_master_awprot;                         // hps_0:h2f_lw_AWPROT -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awprot
	wire  [31:0] hps_0_h2f_lw_axi_master_wdata;                          // hps_0:h2f_lw_WDATA -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wdata
	wire         hps_0_h2f_lw_axi_master_arvalid;                        // hps_0:h2f_lw_ARVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arvalid
	wire   [3:0] hps_0_h2f_lw_axi_master_awcache;                        // hps_0:h2f_lw_AWCACHE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awcache
	wire  [11:0] hps_0_h2f_lw_axi_master_arid;                           // hps_0:h2f_lw_ARID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arid
	wire   [1:0] hps_0_h2f_lw_axi_master_arlock;                         // hps_0:h2f_lw_ARLOCK -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arlock
	wire   [1:0] hps_0_h2f_lw_axi_master_awlock;                         // hps_0:h2f_lw_AWLOCK -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awlock
	wire  [20:0] hps_0_h2f_lw_axi_master_awaddr;                         // hps_0:h2f_lw_AWADDR -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awaddr
	wire   [1:0] hps_0_h2f_lw_axi_master_bresp;                          // mm_interconnect_1:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire         hps_0_h2f_lw_axi_master_arready;                        // mm_interconnect_1:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire  [31:0] hps_0_h2f_lw_axi_master_rdata;                          // mm_interconnect_1:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire         hps_0_h2f_lw_axi_master_awready;                        // mm_interconnect_1:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire   [1:0] hps_0_h2f_lw_axi_master_arburst;                        // hps_0:h2f_lw_ARBURST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arburst
	wire   [2:0] hps_0_h2f_lw_axi_master_arsize;                         // hps_0:h2f_lw_ARSIZE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arsize
	wire         hps_0_h2f_lw_axi_master_bready;                         // hps_0:h2f_lw_BREADY -> mm_interconnect_1:hps_0_h2f_lw_axi_master_bready
	wire         hps_0_h2f_lw_axi_master_rlast;                          // mm_interconnect_1:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire         hps_0_h2f_lw_axi_master_wlast;                          // hps_0:h2f_lw_WLAST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wlast
	wire   [1:0] hps_0_h2f_lw_axi_master_rresp;                          // mm_interconnect_1:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire  [11:0] hps_0_h2f_lw_axi_master_awid;                           // hps_0:h2f_lw_AWID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awid
	wire  [11:0] hps_0_h2f_lw_axi_master_bid;                            // mm_interconnect_1:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire         hps_0_h2f_lw_axi_master_bvalid;                         // mm_interconnect_1:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire   [2:0] hps_0_h2f_lw_axi_master_awsize;                         // hps_0:h2f_lw_AWSIZE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awsize
	wire         hps_0_h2f_lw_axi_master_awvalid;                        // hps_0:h2f_lw_AWVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awvalid
	wire         hps_0_h2f_lw_axi_master_rvalid;                         // mm_interconnect_1:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire         mm_interconnect_1_vga_ball_0_avalon_slave_0_chipselect; // mm_interconnect_1:vga_ball_0_avalon_slave_0_chipselect -> vga_ball_0:chipselect
	wire   [2:0] mm_interconnect_1_vga_ball_0_avalon_slave_0_address;    // mm_interconnect_1:vga_ball_0_avalon_slave_0_address -> vga_ball_0:address
	wire         mm_interconnect_1_vga_ball_0_avalon_slave_0_write;      // mm_interconnect_1:vga_ball_0_avalon_slave_0_write -> vga_ball_0:write
	wire   [7:0] mm_interconnect_1_vga_ball_0_avalon_slave_0_writedata;  // mm_interconnect_1:vga_ball_0_avalon_slave_0_writedata -> vga_ball_0:writedata
	wire  [31:0] hps_0_f2h_irq0_irq;                                     // irq_mapper:sender_irq -> hps_0:f2h_irq_p0
	wire  [31:0] hps_0_f2h_irq1_irq;                                     // irq_mapper_001:sender_irq -> hps_0:f2h_irq_p1
	wire         rst_controller_reset_out_reset;                         // rst_controller:reset_out -> [apple_sprite:reset, map1_0:reset, map1_1:reset, mm_interconnect_0:snake_tail_up_sprite_reset1_reset_bridge_in_reset_reset, mm_interconnect_1:vga_ball_0_reset_reset_bridge_in_reset_reset, rst_translator:in_reset, snake_body_bottomleft_sprite:reset, snake_body_bottomright_sprite:reset, snake_body_horizontal_sprite:reset, snake_body_topleft_sprite:reset, snake_body_topright_sprite:reset, snake_body_vertical_sprite:reset, snake_head_down_sprite:reset, snake_head_left_sprite:reset, snake_head_right_sprite:reset, snake_head_up_sprite:reset, snake_tail_down_sprite:reset, snake_tail_left_sprite:reset, snake_tail_right_sprite:reset, snake_tail_up_sprite:reset, vga_ball_0:reset, wall_sprite:reset]
	wire         rst_controller_reset_out_reset_req;                     // rst_controller:reset_req -> [apple_sprite:reset_req, rst_translator:reset_req_in, snake_body_bottomleft_sprite:reset_req, snake_body_bottomright_sprite:reset_req, snake_body_horizontal_sprite:reset_req, snake_body_topleft_sprite:reset_req, snake_body_topright_sprite:reset_req, snake_body_vertical_sprite:reset_req, snake_head_down_sprite:reset_req, snake_head_left_sprite:reset_req, snake_head_right_sprite:reset_req, snake_head_up_sprite:reset_req, snake_tail_down_sprite:reset_req, snake_tail_left_sprite:reset_req, snake_tail_right_sprite:reset_req, snake_tail_up_sprite:reset_req, wall_sprite:reset_req]
	wire         rst_controller_001_reset_out_reset;                     // rst_controller_001:reset_out -> [mm_interconnect_0:hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset]
	wire         hps_0_h2f_reset_reset;                                  // hps_0:h2f_rst_n -> rst_controller_001:reset_in0

	soc_system_apple_sprite apple_sprite (
		.clk         (clk_clk),                            //   clk1.clk
		.address     (apple_sprite_s1_address),            //     s1.address
		.debugaccess (apple_sprite_s1_debugaccess),        //       .debugaccess
		.clken       (apple_sprite_s1_clken),              //       .clken
		.chipselect  (apple_sprite_s1_chipselect),         //       .chipselect
		.write       (apple_sprite_s1_write),              //       .write
		.readdata    (apple_sprite_s1_readdata),           //       .readdata
		.writedata   (apple_sprite_s1_writedata),          //       .writedata
		.byteenable  (apple_sprite_s1_byteenable),         //       .byteenable
		.reset       (rst_controller_reset_out_reset),     // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req), //       .reset_req
		.freeze      (1'b0)                                // (terminated)
	);

	soc_system_hps_0 #(
		.F2S_Width (2),
		.S2F_Width (2)
	) hps_0 (
		.h2f_user1_clk            (),                                //   h2f_user1_clock.clk
		.mem_a                    (hps_ddr3_mem_a),                  //            memory.mem_a
		.mem_ba                   (hps_ddr3_mem_ba),                 //                  .mem_ba
		.mem_ck                   (hps_ddr3_mem_ck),                 //                  .mem_ck
		.mem_ck_n                 (hps_ddr3_mem_ck_n),               //                  .mem_ck_n
		.mem_cke                  (hps_ddr3_mem_cke),                //                  .mem_cke
		.mem_cs_n                 (hps_ddr3_mem_cs_n),               //                  .mem_cs_n
		.mem_ras_n                (hps_ddr3_mem_ras_n),              //                  .mem_ras_n
		.mem_cas_n                (hps_ddr3_mem_cas_n),              //                  .mem_cas_n
		.mem_we_n                 (hps_ddr3_mem_we_n),               //                  .mem_we_n
		.mem_reset_n              (hps_ddr3_mem_reset_n),            //                  .mem_reset_n
		.mem_dq                   (hps_ddr3_mem_dq),                 //                  .mem_dq
		.mem_dqs                  (hps_ddr3_mem_dqs),                //                  .mem_dqs
		.mem_dqs_n                (hps_ddr3_mem_dqs_n),              //                  .mem_dqs_n
		.mem_odt                  (hps_ddr3_mem_odt),                //                  .mem_odt
		.mem_dm                   (hps_ddr3_mem_dm),                 //                  .mem_dm
		.oct_rzqin                (hps_ddr3_oct_rzqin),              //                  .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_hps_io_emac1_inst_TX_CLK),    //            hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_hps_io_emac1_inst_TXD0),      //                  .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_hps_io_emac1_inst_TXD1),      //                  .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_hps_io_emac1_inst_TXD2),      //                  .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_hps_io_emac1_inst_TXD3),      //                  .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_hps_io_emac1_inst_RXD0),      //                  .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_hps_io_emac1_inst_MDIO),      //                  .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_hps_io_emac1_inst_MDC),       //                  .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_hps_io_emac1_inst_RX_CTL),    //                  .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_hps_io_emac1_inst_TX_CTL),    //                  .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_hps_io_emac1_inst_RX_CLK),    //                  .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_hps_io_emac1_inst_RXD1),      //                  .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_hps_io_emac1_inst_RXD2),      //                  .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_hps_io_emac1_inst_RXD3),      //                  .hps_io_emac1_inst_RXD3
		.hps_io_sdio_inst_CMD     (hps_hps_io_sdio_inst_CMD),        //                  .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_hps_io_sdio_inst_D0),         //                  .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_hps_io_sdio_inst_D1),         //                  .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_hps_io_sdio_inst_CLK),        //                  .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_hps_io_sdio_inst_D2),         //                  .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_hps_io_sdio_inst_D3),         //                  .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_hps_io_usb1_inst_D0),         //                  .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_hps_io_usb1_inst_D1),         //                  .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_hps_io_usb1_inst_D2),         //                  .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_hps_io_usb1_inst_D3),         //                  .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_hps_io_usb1_inst_D4),         //                  .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_hps_io_usb1_inst_D5),         //                  .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_hps_io_usb1_inst_D6),         //                  .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_hps_io_usb1_inst_D7),         //                  .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_hps_io_usb1_inst_CLK),        //                  .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_hps_io_usb1_inst_STP),        //                  .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_hps_io_usb1_inst_DIR),        //                  .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_hps_io_usb1_inst_NXT),        //                  .hps_io_usb1_inst_NXT
		.hps_io_spim1_inst_CLK    (hps_hps_io_spim1_inst_CLK),       //                  .hps_io_spim1_inst_CLK
		.hps_io_spim1_inst_MOSI   (hps_hps_io_spim1_inst_MOSI),      //                  .hps_io_spim1_inst_MOSI
		.hps_io_spim1_inst_MISO   (hps_hps_io_spim1_inst_MISO),      //                  .hps_io_spim1_inst_MISO
		.hps_io_spim1_inst_SS0    (hps_hps_io_spim1_inst_SS0),       //                  .hps_io_spim1_inst_SS0
		.hps_io_uart0_inst_RX     (hps_hps_io_uart0_inst_RX),        //                  .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_hps_io_uart0_inst_TX),        //                  .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_hps_io_i2c0_inst_SDA),        //                  .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_hps_io_i2c0_inst_SCL),        //                  .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA     (hps_hps_io_i2c1_inst_SDA),        //                  .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL     (hps_hps_io_i2c1_inst_SCL),        //                  .hps_io_i2c1_inst_SCL
		.hps_io_gpio_inst_GPIO09  (hps_hps_io_gpio_inst_GPIO09),     //                  .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35  (hps_hps_io_gpio_inst_GPIO35),     //                  .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO40  (hps_hps_io_gpio_inst_GPIO40),     //                  .hps_io_gpio_inst_GPIO40
		.hps_io_gpio_inst_GPIO48  (hps_hps_io_gpio_inst_GPIO48),     //                  .hps_io_gpio_inst_GPIO48
		.hps_io_gpio_inst_GPIO53  (hps_hps_io_gpio_inst_GPIO53),     //                  .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54  (hps_hps_io_gpio_inst_GPIO54),     //                  .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_GPIO61  (hps_hps_io_gpio_inst_GPIO61),     //                  .hps_io_gpio_inst_GPIO61
		.h2f_rst_n                (hps_0_h2f_reset_reset),           //         h2f_reset.reset_n
		.h2f_axi_clk              (clk_clk),                         //     h2f_axi_clock.clk
		.h2f_AWID                 (hps_0_h2f_axi_master_awid),       //    h2f_axi_master.awid
		.h2f_AWADDR               (hps_0_h2f_axi_master_awaddr),     //                  .awaddr
		.h2f_AWLEN                (hps_0_h2f_axi_master_awlen),      //                  .awlen
		.h2f_AWSIZE               (hps_0_h2f_axi_master_awsize),     //                  .awsize
		.h2f_AWBURST              (hps_0_h2f_axi_master_awburst),    //                  .awburst
		.h2f_AWLOCK               (hps_0_h2f_axi_master_awlock),     //                  .awlock
		.h2f_AWCACHE              (hps_0_h2f_axi_master_awcache),    //                  .awcache
		.h2f_AWPROT               (hps_0_h2f_axi_master_awprot),     //                  .awprot
		.h2f_AWVALID              (hps_0_h2f_axi_master_awvalid),    //                  .awvalid
		.h2f_AWREADY              (hps_0_h2f_axi_master_awready),    //                  .awready
		.h2f_WID                  (hps_0_h2f_axi_master_wid),        //                  .wid
		.h2f_WDATA                (hps_0_h2f_axi_master_wdata),      //                  .wdata
		.h2f_WSTRB                (hps_0_h2f_axi_master_wstrb),      //                  .wstrb
		.h2f_WLAST                (hps_0_h2f_axi_master_wlast),      //                  .wlast
		.h2f_WVALID               (hps_0_h2f_axi_master_wvalid),     //                  .wvalid
		.h2f_WREADY               (hps_0_h2f_axi_master_wready),     //                  .wready
		.h2f_BID                  (hps_0_h2f_axi_master_bid),        //                  .bid
		.h2f_BRESP                (hps_0_h2f_axi_master_bresp),      //                  .bresp
		.h2f_BVALID               (hps_0_h2f_axi_master_bvalid),     //                  .bvalid
		.h2f_BREADY               (hps_0_h2f_axi_master_bready),     //                  .bready
		.h2f_ARID                 (hps_0_h2f_axi_master_arid),       //                  .arid
		.h2f_ARADDR               (hps_0_h2f_axi_master_araddr),     //                  .araddr
		.h2f_ARLEN                (hps_0_h2f_axi_master_arlen),      //                  .arlen
		.h2f_ARSIZE               (hps_0_h2f_axi_master_arsize),     //                  .arsize
		.h2f_ARBURST              (hps_0_h2f_axi_master_arburst),    //                  .arburst
		.h2f_ARLOCK               (hps_0_h2f_axi_master_arlock),     //                  .arlock
		.h2f_ARCACHE              (hps_0_h2f_axi_master_arcache),    //                  .arcache
		.h2f_ARPROT               (hps_0_h2f_axi_master_arprot),     //                  .arprot
		.h2f_ARVALID              (hps_0_h2f_axi_master_arvalid),    //                  .arvalid
		.h2f_ARREADY              (hps_0_h2f_axi_master_arready),    //                  .arready
		.h2f_RID                  (hps_0_h2f_axi_master_rid),        //                  .rid
		.h2f_RDATA                (hps_0_h2f_axi_master_rdata),      //                  .rdata
		.h2f_RRESP                (hps_0_h2f_axi_master_rresp),      //                  .rresp
		.h2f_RLAST                (hps_0_h2f_axi_master_rlast),      //                  .rlast
		.h2f_RVALID               (hps_0_h2f_axi_master_rvalid),     //                  .rvalid
		.h2f_RREADY               (hps_0_h2f_axi_master_rready),     //                  .rready
		.f2h_axi_clk              (clk_clk),                         //     f2h_axi_clock.clk
		.f2h_AWID                 (),                                //     f2h_axi_slave.awid
		.f2h_AWADDR               (),                                //                  .awaddr
		.f2h_AWLEN                (),                                //                  .awlen
		.f2h_AWSIZE               (),                                //                  .awsize
		.f2h_AWBURST              (),                                //                  .awburst
		.f2h_AWLOCK               (),                                //                  .awlock
		.f2h_AWCACHE              (),                                //                  .awcache
		.f2h_AWPROT               (),                                //                  .awprot
		.f2h_AWVALID              (),                                //                  .awvalid
		.f2h_AWREADY              (),                                //                  .awready
		.f2h_AWUSER               (),                                //                  .awuser
		.f2h_WID                  (),                                //                  .wid
		.f2h_WDATA                (),                                //                  .wdata
		.f2h_WSTRB                (),                                //                  .wstrb
		.f2h_WLAST                (),                                //                  .wlast
		.f2h_WVALID               (),                                //                  .wvalid
		.f2h_WREADY               (),                                //                  .wready
		.f2h_BID                  (),                                //                  .bid
		.f2h_BRESP                (),                                //                  .bresp
		.f2h_BVALID               (),                                //                  .bvalid
		.f2h_BREADY               (),                                //                  .bready
		.f2h_ARID                 (),                                //                  .arid
		.f2h_ARADDR               (),                                //                  .araddr
		.f2h_ARLEN                (),                                //                  .arlen
		.f2h_ARSIZE               (),                                //                  .arsize
		.f2h_ARBURST              (),                                //                  .arburst
		.f2h_ARLOCK               (),                                //                  .arlock
		.f2h_ARCACHE              (),                                //                  .arcache
		.f2h_ARPROT               (),                                //                  .arprot
		.f2h_ARVALID              (),                                //                  .arvalid
		.f2h_ARREADY              (),                                //                  .arready
		.f2h_ARUSER               (),                                //                  .aruser
		.f2h_RID                  (),                                //                  .rid
		.f2h_RDATA                (),                                //                  .rdata
		.f2h_RRESP                (),                                //                  .rresp
		.f2h_RLAST                (),                                //                  .rlast
		.f2h_RVALID               (),                                //                  .rvalid
		.f2h_RREADY               (),                                //                  .rready
		.h2f_lw_axi_clk           (clk_clk),                         //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (hps_0_h2f_lw_axi_master_awid),    // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (hps_0_h2f_lw_axi_master_awaddr),  //                  .awaddr
		.h2f_lw_AWLEN             (hps_0_h2f_lw_axi_master_awlen),   //                  .awlen
		.h2f_lw_AWSIZE            (hps_0_h2f_lw_axi_master_awsize),  //                  .awsize
		.h2f_lw_AWBURST           (hps_0_h2f_lw_axi_master_awburst), //                  .awburst
		.h2f_lw_AWLOCK            (hps_0_h2f_lw_axi_master_awlock),  //                  .awlock
		.h2f_lw_AWCACHE           (hps_0_h2f_lw_axi_master_awcache), //                  .awcache
		.h2f_lw_AWPROT            (hps_0_h2f_lw_axi_master_awprot),  //                  .awprot
		.h2f_lw_AWVALID           (hps_0_h2f_lw_axi_master_awvalid), //                  .awvalid
		.h2f_lw_AWREADY           (hps_0_h2f_lw_axi_master_awready), //                  .awready
		.h2f_lw_WID               (hps_0_h2f_lw_axi_master_wid),     //                  .wid
		.h2f_lw_WDATA             (hps_0_h2f_lw_axi_master_wdata),   //                  .wdata
		.h2f_lw_WSTRB             (hps_0_h2f_lw_axi_master_wstrb),   //                  .wstrb
		.h2f_lw_WLAST             (hps_0_h2f_lw_axi_master_wlast),   //                  .wlast
		.h2f_lw_WVALID            (hps_0_h2f_lw_axi_master_wvalid),  //                  .wvalid
		.h2f_lw_WREADY            (hps_0_h2f_lw_axi_master_wready),  //                  .wready
		.h2f_lw_BID               (hps_0_h2f_lw_axi_master_bid),     //                  .bid
		.h2f_lw_BRESP             (hps_0_h2f_lw_axi_master_bresp),   //                  .bresp
		.h2f_lw_BVALID            (hps_0_h2f_lw_axi_master_bvalid),  //                  .bvalid
		.h2f_lw_BREADY            (hps_0_h2f_lw_axi_master_bready),  //                  .bready
		.h2f_lw_ARID              (hps_0_h2f_lw_axi_master_arid),    //                  .arid
		.h2f_lw_ARADDR            (hps_0_h2f_lw_axi_master_araddr),  //                  .araddr
		.h2f_lw_ARLEN             (hps_0_h2f_lw_axi_master_arlen),   //                  .arlen
		.h2f_lw_ARSIZE            (hps_0_h2f_lw_axi_master_arsize),  //                  .arsize
		.h2f_lw_ARBURST           (hps_0_h2f_lw_axi_master_arburst), //                  .arburst
		.h2f_lw_ARLOCK            (hps_0_h2f_lw_axi_master_arlock),  //                  .arlock
		.h2f_lw_ARCACHE           (hps_0_h2f_lw_axi_master_arcache), //                  .arcache
		.h2f_lw_ARPROT            (hps_0_h2f_lw_axi_master_arprot),  //                  .arprot
		.h2f_lw_ARVALID           (hps_0_h2f_lw_axi_master_arvalid), //                  .arvalid
		.h2f_lw_ARREADY           (hps_0_h2f_lw_axi_master_arready), //                  .arready
		.h2f_lw_RID               (hps_0_h2f_lw_axi_master_rid),     //                  .rid
		.h2f_lw_RDATA             (hps_0_h2f_lw_axi_master_rdata),   //                  .rdata
		.h2f_lw_RRESP             (hps_0_h2f_lw_axi_master_rresp),   //                  .rresp
		.h2f_lw_RLAST             (hps_0_h2f_lw_axi_master_rlast),   //                  .rlast
		.h2f_lw_RVALID            (hps_0_h2f_lw_axi_master_rvalid),  //                  .rvalid
		.h2f_lw_RREADY            (hps_0_h2f_lw_axi_master_rready),  //                  .rready
		.f2h_irq_p0               (hps_0_f2h_irq0_irq),              //          f2h_irq0.irq
		.f2h_irq_p1               (hps_0_f2h_irq1_irq)               //          f2h_irq1.irq
	);

	vga_ball map1_0 (
		.clk         (clk_clk),                          //          clock.clk
		.reset       (rst_controller_reset_out_reset),   //          reset.reset
		.address     (map1_0_avalon_slave_0_address),    // avalon_slave_0.address
		.chipselect  (map1_0_avalon_slave_0_chipselect), //               .chipselect
		.write       (map1_0_avalon_slave_0_write),      //               .write
		.writedata   (map1_0_avalon_slave_0_writedata),  //               .writedata
		.VGA_B       (map1_0_vga_b),                     //            vga.b
		.VGA_BLANK_n (map1_0_vga_blank_n),               //               .blank_n
		.VGA_CLK     (map1_0_vga_clk),                   //               .clk
		.VGA_G       (map1_0_vga_g),                     //               .g
		.VGA_HS      (map1_0_vga_hs),                    //               .hs
		.VGA_R       (map1_0_vga_r),                     //               .r
		.VGA_SYNC_n  (map1_0_vga_sync_n),                //               .sync_n
		.VGA_VS      (map1_0_vga_vs)                     //               .vs
	);

	vga_ball map1_1 (
		.clk         (clk_clk),                          //          clock.clk
		.reset       (rst_controller_reset_out_reset),   //          reset.reset
		.address     (map1_1_avalon_slave_0_address),    // avalon_slave_0.address
		.chipselect  (map1_1_avalon_slave_0_chipselect), //               .chipselect
		.write       (map1_1_avalon_slave_0_write),      //               .write
		.writedata   (map1_1_avalon_slave_0_writedata),  //               .writedata
		.VGA_B       (map1_1_vga_b),                     //            vga.b
		.VGA_BLANK_n (map1_1_vga_blank_n),               //               .blank_n
		.VGA_CLK     (map1_1_vga_clk),                   //               .clk
		.VGA_G       (map1_1_vga_g),                     //               .g
		.VGA_HS      (map1_1_vga_hs),                    //               .hs
		.VGA_R       (map1_1_vga_r),                     //               .r
		.VGA_SYNC_n  (map1_1_vga_sync_n),                //               .sync_n
		.VGA_VS      (map1_1_vga_vs)                     //               .vs
	);

	soc_system_snake_body_bottomleft_sprite snake_body_bottomleft_sprite (
		.clk         (clk_clk),                                     //   clk1.clk
		.address     (snake_body_bottomleft_sprite_s1_address),     //     s1.address
		.debugaccess (snake_body_bottomleft_sprite_s1_debugaccess), //       .debugaccess
		.clken       (snake_body_bottomleft_sprite_s1_clken),       //       .clken
		.chipselect  (snake_body_bottomleft_sprite_s1_chipselect),  //       .chipselect
		.write       (snake_body_bottomleft_sprite_s1_write),       //       .write
		.readdata    (snake_body_bottomleft_sprite_s1_readdata),    //       .readdata
		.writedata   (snake_body_bottomleft_sprite_s1_writedata),   //       .writedata
		.byteenable  (snake_body_bottomleft_sprite_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),              // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),          //       .reset_req
		.freeze      (1'b0)                                         // (terminated)
	);

	soc_system_snake_body_bottomright_sprite snake_body_bottomright_sprite (
		.clk         (clk_clk),                                      //   clk1.clk
		.address     (snake_body_bottomright_sprite_s1_address),     //     s1.address
		.debugaccess (snake_body_bottomright_sprite_s1_debugaccess), //       .debugaccess
		.clken       (snake_body_bottomright_sprite_s1_clken),       //       .clken
		.chipselect  (snake_body_bottomright_sprite_s1_chipselect),  //       .chipselect
		.write       (snake_body_bottomright_sprite_s1_write),       //       .write
		.readdata    (snake_body_bottomright_sprite_s1_readdata),    //       .readdata
		.writedata   (snake_body_bottomright_sprite_s1_writedata),   //       .writedata
		.byteenable  (snake_body_bottomright_sprite_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),               // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),           //       .reset_req
		.freeze      (1'b0)                                          // (terminated)
	);

	soc_system_snake_body_horizontal_sprite snake_body_horizontal_sprite (
		.clk         (clk_clk),                                     //   clk1.clk
		.address     (snake_body_horizontal_sprite_s1_address),     //     s1.address
		.debugaccess (snake_body_horizontal_sprite_s1_debugaccess), //       .debugaccess
		.clken       (snake_body_horizontal_sprite_s1_clken),       //       .clken
		.chipselect  (snake_body_horizontal_sprite_s1_chipselect),  //       .chipselect
		.write       (snake_body_horizontal_sprite_s1_write),       //       .write
		.readdata    (snake_body_horizontal_sprite_s1_readdata),    //       .readdata
		.writedata   (snake_body_horizontal_sprite_s1_writedata),   //       .writedata
		.byteenable  (snake_body_horizontal_sprite_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),              // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),          //       .reset_req
		.freeze      (1'b0)                                         // (terminated)
	);

	soc_system_snake_body_topleft_sprite snake_body_topleft_sprite (
		.clk         (clk_clk),                                  //   clk1.clk
		.address     (snake_body_topleft_sprite_s1_address),     //     s1.address
		.debugaccess (snake_body_topleft_sprite_s1_debugaccess), //       .debugaccess
		.clken       (snake_body_topleft_sprite_s1_clken),       //       .clken
		.chipselect  (snake_body_topleft_sprite_s1_chipselect),  //       .chipselect
		.write       (snake_body_topleft_sprite_s1_write),       //       .write
		.readdata    (snake_body_topleft_sprite_s1_readdata),    //       .readdata
		.writedata   (snake_body_topleft_sprite_s1_writedata),   //       .writedata
		.byteenable  (snake_body_topleft_sprite_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),           // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),       //       .reset_req
		.freeze      (1'b0)                                      // (terminated)
	);

	soc_system_snake_body_topright_sprite snake_body_topright_sprite (
		.clk         (clk_clk),                                   //   clk1.clk
		.address     (snake_body_topright_sprite_s1_address),     //     s1.address
		.debugaccess (snake_body_topright_sprite_s1_debugaccess), //       .debugaccess
		.clken       (snake_body_topright_sprite_s1_clken),       //       .clken
		.chipselect  (snake_body_topright_sprite_s1_chipselect),  //       .chipselect
		.write       (snake_body_topright_sprite_s1_write),       //       .write
		.readdata    (snake_body_topright_sprite_s1_readdata),    //       .readdata
		.writedata   (snake_body_topright_sprite_s1_writedata),   //       .writedata
		.byteenable  (snake_body_topright_sprite_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),            // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),        //       .reset_req
		.freeze      (1'b0)                                       // (terminated)
	);

	soc_system_snake_body_vertical_sprite snake_body_vertical_sprite (
		.clk         (clk_clk),                                   //   clk1.clk
		.address     (snake_body_vertical_sprite_s1_address),     //     s1.address
		.debugaccess (snake_body_vertical_sprite_s1_debugaccess), //       .debugaccess
		.clken       (snake_body_vertical_sprite_s1_clken),       //       .clken
		.chipselect  (snake_body_vertical_sprite_s1_chipselect),  //       .chipselect
		.write       (snake_body_vertical_sprite_s1_write),       //       .write
		.readdata    (snake_body_vertical_sprite_s1_readdata),    //       .readdata
		.writedata   (snake_body_vertical_sprite_s1_writedata),   //       .writedata
		.byteenable  (snake_body_vertical_sprite_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),            // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),        //       .reset_req
		.freeze      (1'b0)                                       // (terminated)
	);

	soc_system_snake_head_down_sprite snake_head_down_sprite (
		.clk         (clk_clk),                               //   clk1.clk
		.address     (snake_head_down_sprite_s1_address),     //     s1.address
		.debugaccess (snake_head_down_sprite_s1_debugaccess), //       .debugaccess
		.clken       (snake_head_down_sprite_s1_clken),       //       .clken
		.chipselect  (snake_head_down_sprite_s1_chipselect),  //       .chipselect
		.write       (snake_head_down_sprite_s1_write),       //       .write
		.readdata    (snake_head_down_sprite_s1_readdata),    //       .readdata
		.writedata   (snake_head_down_sprite_s1_writedata),   //       .writedata
		.byteenable  (snake_head_down_sprite_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),        // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),    //       .reset_req
		.freeze      (1'b0)                                   // (terminated)
	);

	soc_system_snake_head_left_sprite snake_head_left_sprite (
		.clk         (clk_clk),                               //   clk1.clk
		.address     (snake_head_left_sprite_s1_address),     //     s1.address
		.debugaccess (snake_head_left_sprite_s1_debugaccess), //       .debugaccess
		.clken       (snake_head_left_sprite_s1_clken),       //       .clken
		.chipselect  (snake_head_left_sprite_s1_chipselect),  //       .chipselect
		.write       (snake_head_left_sprite_s1_write),       //       .write
		.readdata    (snake_head_left_sprite_s1_readdata),    //       .readdata
		.writedata   (snake_head_left_sprite_s1_writedata),   //       .writedata
		.byteenable  (snake_head_left_sprite_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),        // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),    //       .reset_req
		.freeze      (1'b0)                                   // (terminated)
	);

	soc_system_snake_head_right_sprite snake_head_right_sprite (
		.clk         (clk_clk),                                //   clk1.clk
		.address     (snake_head_right_sprite_s1_address),     //     s1.address
		.debugaccess (snake_head_right_sprite_s1_debugaccess), //       .debugaccess
		.clken       (snake_head_right_sprite_s1_clken),       //       .clken
		.chipselect  (snake_head_right_sprite_s1_chipselect),  //       .chipselect
		.write       (snake_head_right_sprite_s1_write),       //       .write
		.readdata    (snake_head_right_sprite_s1_readdata),    //       .readdata
		.writedata   (snake_head_right_sprite_s1_writedata),   //       .writedata
		.byteenable  (snake_head_right_sprite_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),         // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),     //       .reset_req
		.freeze      (1'b0)                                    // (terminated)
	);

	soc_system_snake_head_up_sprite snake_head_up_sprite (
		.clk         (clk_clk),                             //   clk1.clk
		.address     (snake_head_up_sprite_s1_address),     //     s1.address
		.debugaccess (snake_head_up_sprite_s1_debugaccess), //       .debugaccess
		.clken       (snake_head_up_sprite_s1_clken),       //       .clken
		.chipselect  (snake_head_up_sprite_s1_chipselect),  //       .chipselect
		.write       (snake_head_up_sprite_s1_write),       //       .write
		.readdata    (snake_head_up_sprite_s1_readdata),    //       .readdata
		.writedata   (snake_head_up_sprite_s1_writedata),   //       .writedata
		.byteenable  (snake_head_up_sprite_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),  //       .reset_req
		.freeze      (1'b0)                                 // (terminated)
	);

	soc_system_snake_tail_down_sprite snake_tail_down_sprite (
		.clk         (clk_clk),                               //   clk1.clk
		.address     (snake_tail_down_sprite_s1_address),     //     s1.address
		.debugaccess (snake_tail_down_sprite_s1_debugaccess), //       .debugaccess
		.clken       (snake_tail_down_sprite_s1_clken),       //       .clken
		.chipselect  (snake_tail_down_sprite_s1_chipselect),  //       .chipselect
		.write       (snake_tail_down_sprite_s1_write),       //       .write
		.readdata    (snake_tail_down_sprite_s1_readdata),    //       .readdata
		.writedata   (snake_tail_down_sprite_s1_writedata),   //       .writedata
		.byteenable  (snake_tail_down_sprite_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),        // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),    //       .reset_req
		.freeze      (1'b0)                                   // (terminated)
	);

	soc_system_snake_tail_left_sprite snake_tail_left_sprite (
		.clk         (clk_clk),                               //   clk1.clk
		.address     (snake_tail_left_sprite_s1_address),     //     s1.address
		.debugaccess (snake_tail_left_sprite_s1_debugaccess), //       .debugaccess
		.clken       (snake_tail_left_sprite_s1_clken),       //       .clken
		.chipselect  (snake_tail_left_sprite_s1_chipselect),  //       .chipselect
		.write       (snake_tail_left_sprite_s1_write),       //       .write
		.readdata    (snake_tail_left_sprite_s1_readdata),    //       .readdata
		.writedata   (snake_tail_left_sprite_s1_writedata),   //       .writedata
		.byteenable  (snake_tail_left_sprite_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),        // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),    //       .reset_req
		.freeze      (1'b0)                                   // (terminated)
	);

	soc_system_snake_tail_right_sprite snake_tail_right_sprite (
		.clk         (clk_clk),                                //   clk1.clk
		.address     (snake_tail_right_sprite_s1_address),     //     s1.address
		.debugaccess (snake_tail_right_sprite_s1_debugaccess), //       .debugaccess
		.clken       (snake_tail_right_sprite_s1_clken),       //       .clken
		.chipselect  (snake_tail_right_sprite_s1_chipselect),  //       .chipselect
		.write       (snake_tail_right_sprite_s1_write),       //       .write
		.readdata    (snake_tail_right_sprite_s1_readdata),    //       .readdata
		.writedata   (snake_tail_right_sprite_s1_writedata),   //       .writedata
		.byteenable  (snake_tail_right_sprite_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),         // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),     //       .reset_req
		.freeze      (1'b0)                                    // (terminated)
	);

	soc_system_snake_tail_up_sprite snake_tail_up_sprite (
		.clk         (clk_clk),                                               //   clk1.clk
		.address     (mm_interconnect_0_snake_tail_up_sprite_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_snake_tail_up_sprite_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_snake_tail_up_sprite_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_snake_tail_up_sprite_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_snake_tail_up_sprite_s1_write),       //       .write
		.readdata    (mm_interconnect_0_snake_tail_up_sprite_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_snake_tail_up_sprite_s1_writedata),   //       .writedata
		.byteenable  (mm_interconnect_0_snake_tail_up_sprite_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),                        // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),                    //       .reset_req
		.freeze      (1'b0)                                                   // (terminated)
	);

	vga_ball vga_ball_0 (
		.clk         (clk_clk),                                                //          clock.clk
		.reset       (rst_controller_reset_out_reset),                         //          reset.reset
		.VGA_B       (vga_b),                                                  //            vga.b
		.VGA_BLANK_n (vga_blank_n),                                            //               .blank_n
		.VGA_CLK     (vga_clk),                                                //               .clk
		.VGA_G       (vga_g),                                                  //               .g
		.VGA_HS      (vga_hs),                                                 //               .hs
		.VGA_R       (vga_r),                                                  //               .r
		.VGA_SYNC_n  (vga_sync_n),                                             //               .sync_n
		.VGA_VS      (vga_vs),                                                 //               .vs
		.writedata   (mm_interconnect_1_vga_ball_0_avalon_slave_0_writedata),  // avalon_slave_0.writedata
		.write       (mm_interconnect_1_vga_ball_0_avalon_slave_0_write),      //               .write
		.chipselect  (mm_interconnect_1_vga_ball_0_avalon_slave_0_chipselect), //               .chipselect
		.address     (mm_interconnect_1_vga_ball_0_avalon_slave_0_address)     //               .address
	);

	soc_system_wall_sprite wall_sprite (
		.clk         (clk_clk),                            //   clk1.clk
		.address     (wall_sprite_s1_address),             //     s1.address
		.debugaccess (wall_sprite_s1_debugaccess),         //       .debugaccess
		.clken       (wall_sprite_s1_clken),               //       .clken
		.chipselect  (wall_sprite_s1_chipselect),          //       .chipselect
		.write       (wall_sprite_s1_write),               //       .write
		.readdata    (wall_sprite_s1_readdata),            //       .readdata
		.writedata   (wall_sprite_s1_writedata),           //       .writedata
		.byteenable  (wall_sprite_s1_byteenable),          //       .byteenable
		.reset       (rst_controller_reset_out_reset),     // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req), //       .reset_req
		.freeze      (1'b0)                                // (terminated)
	);

	soc_system_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_h2f_axi_master_awid                                        (hps_0_h2f_axi_master_awid),                             //                                       hps_0_h2f_axi_master.awid
		.hps_0_h2f_axi_master_awaddr                                      (hps_0_h2f_axi_master_awaddr),                           //                                                           .awaddr
		.hps_0_h2f_axi_master_awlen                                       (hps_0_h2f_axi_master_awlen),                            //                                                           .awlen
		.hps_0_h2f_axi_master_awsize                                      (hps_0_h2f_axi_master_awsize),                           //                                                           .awsize
		.hps_0_h2f_axi_master_awburst                                     (hps_0_h2f_axi_master_awburst),                          //                                                           .awburst
		.hps_0_h2f_axi_master_awlock                                      (hps_0_h2f_axi_master_awlock),                           //                                                           .awlock
		.hps_0_h2f_axi_master_awcache                                     (hps_0_h2f_axi_master_awcache),                          //                                                           .awcache
		.hps_0_h2f_axi_master_awprot                                      (hps_0_h2f_axi_master_awprot),                           //                                                           .awprot
		.hps_0_h2f_axi_master_awvalid                                     (hps_0_h2f_axi_master_awvalid),                          //                                                           .awvalid
		.hps_0_h2f_axi_master_awready                                     (hps_0_h2f_axi_master_awready),                          //                                                           .awready
		.hps_0_h2f_axi_master_wid                                         (hps_0_h2f_axi_master_wid),                              //                                                           .wid
		.hps_0_h2f_axi_master_wdata                                       (hps_0_h2f_axi_master_wdata),                            //                                                           .wdata
		.hps_0_h2f_axi_master_wstrb                                       (hps_0_h2f_axi_master_wstrb),                            //                                                           .wstrb
		.hps_0_h2f_axi_master_wlast                                       (hps_0_h2f_axi_master_wlast),                            //                                                           .wlast
		.hps_0_h2f_axi_master_wvalid                                      (hps_0_h2f_axi_master_wvalid),                           //                                                           .wvalid
		.hps_0_h2f_axi_master_wready                                      (hps_0_h2f_axi_master_wready),                           //                                                           .wready
		.hps_0_h2f_axi_master_bid                                         (hps_0_h2f_axi_master_bid),                              //                                                           .bid
		.hps_0_h2f_axi_master_bresp                                       (hps_0_h2f_axi_master_bresp),                            //                                                           .bresp
		.hps_0_h2f_axi_master_bvalid                                      (hps_0_h2f_axi_master_bvalid),                           //                                                           .bvalid
		.hps_0_h2f_axi_master_bready                                      (hps_0_h2f_axi_master_bready),                           //                                                           .bready
		.hps_0_h2f_axi_master_arid                                        (hps_0_h2f_axi_master_arid),                             //                                                           .arid
		.hps_0_h2f_axi_master_araddr                                      (hps_0_h2f_axi_master_araddr),                           //                                                           .araddr
		.hps_0_h2f_axi_master_arlen                                       (hps_0_h2f_axi_master_arlen),                            //                                                           .arlen
		.hps_0_h2f_axi_master_arsize                                      (hps_0_h2f_axi_master_arsize),                           //                                                           .arsize
		.hps_0_h2f_axi_master_arburst                                     (hps_0_h2f_axi_master_arburst),                          //                                                           .arburst
		.hps_0_h2f_axi_master_arlock                                      (hps_0_h2f_axi_master_arlock),                           //                                                           .arlock
		.hps_0_h2f_axi_master_arcache                                     (hps_0_h2f_axi_master_arcache),                          //                                                           .arcache
		.hps_0_h2f_axi_master_arprot                                      (hps_0_h2f_axi_master_arprot),                           //                                                           .arprot
		.hps_0_h2f_axi_master_arvalid                                     (hps_0_h2f_axi_master_arvalid),                          //                                                           .arvalid
		.hps_0_h2f_axi_master_arready                                     (hps_0_h2f_axi_master_arready),                          //                                                           .arready
		.hps_0_h2f_axi_master_rid                                         (hps_0_h2f_axi_master_rid),                              //                                                           .rid
		.hps_0_h2f_axi_master_rdata                                       (hps_0_h2f_axi_master_rdata),                            //                                                           .rdata
		.hps_0_h2f_axi_master_rresp                                       (hps_0_h2f_axi_master_rresp),                            //                                                           .rresp
		.hps_0_h2f_axi_master_rlast                                       (hps_0_h2f_axi_master_rlast),                            //                                                           .rlast
		.hps_0_h2f_axi_master_rvalid                                      (hps_0_h2f_axi_master_rvalid),                           //                                                           .rvalid
		.hps_0_h2f_axi_master_rready                                      (hps_0_h2f_axi_master_rready),                           //                                                           .rready
		.clk_0_clk_clk                                                    (clk_clk),                                               //                                                  clk_0_clk.clk
		.hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                    // hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.snake_tail_up_sprite_reset1_reset_bridge_in_reset_reset          (rst_controller_reset_out_reset),                        //          snake_tail_up_sprite_reset1_reset_bridge_in_reset.reset
		.snake_tail_up_sprite_s1_address                                  (mm_interconnect_0_snake_tail_up_sprite_s1_address),     //                                    snake_tail_up_sprite_s1.address
		.snake_tail_up_sprite_s1_write                                    (mm_interconnect_0_snake_tail_up_sprite_s1_write),       //                                                           .write
		.snake_tail_up_sprite_s1_readdata                                 (mm_interconnect_0_snake_tail_up_sprite_s1_readdata),    //                                                           .readdata
		.snake_tail_up_sprite_s1_writedata                                (mm_interconnect_0_snake_tail_up_sprite_s1_writedata),   //                                                           .writedata
		.snake_tail_up_sprite_s1_byteenable                               (mm_interconnect_0_snake_tail_up_sprite_s1_byteenable),  //                                                           .byteenable
		.snake_tail_up_sprite_s1_chipselect                               (mm_interconnect_0_snake_tail_up_sprite_s1_chipselect),  //                                                           .chipselect
		.snake_tail_up_sprite_s1_clken                                    (mm_interconnect_0_snake_tail_up_sprite_s1_clken),       //                                                           .clken
		.snake_tail_up_sprite_s1_debugaccess                              (mm_interconnect_0_snake_tail_up_sprite_s1_debugaccess)  //                                                           .debugaccess
	);

	soc_system_mm_interconnect_1 mm_interconnect_1 (
		.hps_0_h2f_lw_axi_master_awid                                        (hps_0_h2f_lw_axi_master_awid),                           //                                       hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                                      (hps_0_h2f_lw_axi_master_awaddr),                         //                                                              .awaddr
		.hps_0_h2f_lw_axi_master_awlen                                       (hps_0_h2f_lw_axi_master_awlen),                          //                                                              .awlen
		.hps_0_h2f_lw_axi_master_awsize                                      (hps_0_h2f_lw_axi_master_awsize),                         //                                                              .awsize
		.hps_0_h2f_lw_axi_master_awburst                                     (hps_0_h2f_lw_axi_master_awburst),                        //                                                              .awburst
		.hps_0_h2f_lw_axi_master_awlock                                      (hps_0_h2f_lw_axi_master_awlock),                         //                                                              .awlock
		.hps_0_h2f_lw_axi_master_awcache                                     (hps_0_h2f_lw_axi_master_awcache),                        //                                                              .awcache
		.hps_0_h2f_lw_axi_master_awprot                                      (hps_0_h2f_lw_axi_master_awprot),                         //                                                              .awprot
		.hps_0_h2f_lw_axi_master_awvalid                                     (hps_0_h2f_lw_axi_master_awvalid),                        //                                                              .awvalid
		.hps_0_h2f_lw_axi_master_awready                                     (hps_0_h2f_lw_axi_master_awready),                        //                                                              .awready
		.hps_0_h2f_lw_axi_master_wid                                         (hps_0_h2f_lw_axi_master_wid),                            //                                                              .wid
		.hps_0_h2f_lw_axi_master_wdata                                       (hps_0_h2f_lw_axi_master_wdata),                          //                                                              .wdata
		.hps_0_h2f_lw_axi_master_wstrb                                       (hps_0_h2f_lw_axi_master_wstrb),                          //                                                              .wstrb
		.hps_0_h2f_lw_axi_master_wlast                                       (hps_0_h2f_lw_axi_master_wlast),                          //                                                              .wlast
		.hps_0_h2f_lw_axi_master_wvalid                                      (hps_0_h2f_lw_axi_master_wvalid),                         //                                                              .wvalid
		.hps_0_h2f_lw_axi_master_wready                                      (hps_0_h2f_lw_axi_master_wready),                         //                                                              .wready
		.hps_0_h2f_lw_axi_master_bid                                         (hps_0_h2f_lw_axi_master_bid),                            //                                                              .bid
		.hps_0_h2f_lw_axi_master_bresp                                       (hps_0_h2f_lw_axi_master_bresp),                          //                                                              .bresp
		.hps_0_h2f_lw_axi_master_bvalid                                      (hps_0_h2f_lw_axi_master_bvalid),                         //                                                              .bvalid
		.hps_0_h2f_lw_axi_master_bready                                      (hps_0_h2f_lw_axi_master_bready),                         //                                                              .bready
		.hps_0_h2f_lw_axi_master_arid                                        (hps_0_h2f_lw_axi_master_arid),                           //                                                              .arid
		.hps_0_h2f_lw_axi_master_araddr                                      (hps_0_h2f_lw_axi_master_araddr),                         //                                                              .araddr
		.hps_0_h2f_lw_axi_master_arlen                                       (hps_0_h2f_lw_axi_master_arlen),                          //                                                              .arlen
		.hps_0_h2f_lw_axi_master_arsize                                      (hps_0_h2f_lw_axi_master_arsize),                         //                                                              .arsize
		.hps_0_h2f_lw_axi_master_arburst                                     (hps_0_h2f_lw_axi_master_arburst),                        //                                                              .arburst
		.hps_0_h2f_lw_axi_master_arlock                                      (hps_0_h2f_lw_axi_master_arlock),                         //                                                              .arlock
		.hps_0_h2f_lw_axi_master_arcache                                     (hps_0_h2f_lw_axi_master_arcache),                        //                                                              .arcache
		.hps_0_h2f_lw_axi_master_arprot                                      (hps_0_h2f_lw_axi_master_arprot),                         //                                                              .arprot
		.hps_0_h2f_lw_axi_master_arvalid                                     (hps_0_h2f_lw_axi_master_arvalid),                        //                                                              .arvalid
		.hps_0_h2f_lw_axi_master_arready                                     (hps_0_h2f_lw_axi_master_arready),                        //                                                              .arready
		.hps_0_h2f_lw_axi_master_rid                                         (hps_0_h2f_lw_axi_master_rid),                            //                                                              .rid
		.hps_0_h2f_lw_axi_master_rdata                                       (hps_0_h2f_lw_axi_master_rdata),                          //                                                              .rdata
		.hps_0_h2f_lw_axi_master_rresp                                       (hps_0_h2f_lw_axi_master_rresp),                          //                                                              .rresp
		.hps_0_h2f_lw_axi_master_rlast                                       (hps_0_h2f_lw_axi_master_rlast),                          //                                                              .rlast
		.hps_0_h2f_lw_axi_master_rvalid                                      (hps_0_h2f_lw_axi_master_rvalid),                         //                                                              .rvalid
		.hps_0_h2f_lw_axi_master_rready                                      (hps_0_h2f_lw_axi_master_rready),                         //                                                              .rready
		.clk_0_clk_clk                                                       (clk_clk),                                                //                                                     clk_0_clk.clk
		.hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                     // hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.vga_ball_0_reset_reset_bridge_in_reset_reset                        (rst_controller_reset_out_reset),                         //                        vga_ball_0_reset_reset_bridge_in_reset.reset
		.vga_ball_0_avalon_slave_0_address                                   (mm_interconnect_1_vga_ball_0_avalon_slave_0_address),    //                                     vga_ball_0_avalon_slave_0.address
		.vga_ball_0_avalon_slave_0_write                                     (mm_interconnect_1_vga_ball_0_avalon_slave_0_write),      //                                                              .write
		.vga_ball_0_avalon_slave_0_writedata                                 (mm_interconnect_1_vga_ball_0_avalon_slave_0_writedata),  //                                                              .writedata
		.vga_ball_0_avalon_slave_0_chipselect                                (mm_interconnect_1_vga_ball_0_avalon_slave_0_chipselect)  //                                                              .chipselect
	);

	soc_system_irq_mapper irq_mapper (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq0_irq)  //    sender.irq
	);

	soc_system_irq_mapper irq_mapper_001 (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq1_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
